bind async
