`define DSIZE 8
`define ASIZE 4
`define DEPTH 2**`ASIZE
`define no_of_transaction 20
